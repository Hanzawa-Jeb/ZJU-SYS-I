module Mux4T1_32(
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    input [31:0] I3,
    input [1:0] S,
    output [31:0] O
);

Mux4T1_1(I0[0], I1[0], I2[0], I3[0], O[0], S);
Mux4T1_1(I0[1], I1[1], I2[1], I3[1], O[1], S);
Mux4T1_1(I0[2], I1[2], I2[2], I3[2], O[2], S);
Mux4T1_1(I0[3], I1[3], I2[3], I3[3], O[3], S);
Mux4T1_1(I0[4], I1[4], I2[4], I3[4], O[4], S);
Mux4T1_1(I0[5], I1[5], I2[5], I3[5], O[5], S);
Mux4T1_1(I0[6], I1[6], I2[6], I3[6], O[6], S);
Mux4T1_1(I0[7], I1[7], I2[7], I3[7], O[7], S);
Mux4T1_1(I0[8], I1[8], I2[8], I3[8], O[8], S);
Mux4T1_1(I0[9], I1[9], I2[9], I3[9], O[9], S);
Mux4T1_1(I0[10], I1[10], I2[10], I3[10], O[10], S);
Mux4T1_1(I0[11], I1[11], I2[11], I3[11], O[11], S);
Mux4T1_1(I0[12], I1[12], I2[12], I3[12], O[12], S);
Mux4T1_1(I0[13], I1[13], I2[13], I3[13], O[13], S);
Mux4T1_1(I0[14], I1[14], I2[14], I3[14], O[14], S);
Mux4T1_1(I0[15], I1[15], I2[15], I3[15], O[15], S);
Mux4T1_1(I0[16], I1[16], I2[16], I3[16], O[16], S);
Mux4T1_1(I0[17], I1[17], I2[17], I3[17], O[17], S);
Mux4T1_1(I0[18], I1[18], I2[18], I3[18], O[18], S);
Mux4T1_1(I0[19], I1[19], I2[19], I3[19], O[19], S);
Mux4T1_1(I0[20], I1[20], I2[20], I3[20], O[20], S);
Mux4T1_1(I0[21], I1[21], I2[21], I3[21], O[21], S);
Mux4T1_1(I0[22], I1[22], I2[22], I3[22], O[22], S);
Mux4T1_1(I0[23], I1[23], I2[23], I3[23], O[23], S);
Mux4T1_1(I0[24], I1[24], I2[24], I3[24], O[24], S);
Mux4T1_1(I0[25], I1[25], I2[25], I3[25], O[25], S);
Mux4T1_1(I0[26], I1[26], I2[26], I3[26], O[26], S);
Mux4T1_1(I0[27], I1[27], I2[27], I3[27], O[27], S);
Mux4T1_1(I0[28], I1[28], I2[28], I3[28], O[28], S);
Mux4T1_1(I0[29], I1[29], I2[29], I3[29], O[29], S);
Mux4T1_1(I0[30], I1[30], I2[30], I3[30], O[30], S);
Mux4T1_1(I0[31], I1[31], I2[31], I3[31], O[31], S);


    //fill your code

endmodule

